0
0 0 0 0 0 r 68 70 h 1 B 51 B
10 10 10 10 10 r h 6 B 48 B
10 10 10 13 10 r h 11 B 36 B
10 10 10 10 10 r h 23 B 39 B
3 10 0 8 4 8 3 5 3 3 1 6 2 4 5 7 0 4 4 11 1 11 1 3 4 9 3 2 0 10 2 5 2 6 2 12 4 9
-1
